** Profile: "SCHEMATIC1-simulacion_mayor_0.7"  [ D:\TRABAJO ELECTRONICA 19-20\Circuito proteccion\circuito proteccion-pspicefiles\schematic1\simulacion_mayor_0.7.sim ] 

** Creating circuit file "simulacion_mayor_0.7.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Capture_Cis\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
